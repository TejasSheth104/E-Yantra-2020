module TWS(
	input s1, s2,
	output z
);

assign z = (s1^s2);

endmodule
